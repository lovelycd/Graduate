module Four_Vote_74hc151_2_8(input En,A,B,C,D,output F);
	Coder_8_3_74hc151_2_7 C83_151_27_1(En,0,A,B,C,0,D,0,1,0,1,D,1,F);
endmodule 